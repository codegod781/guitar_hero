/*
 * Avalon memory-mapped peripheral that generates VGA
 *
 * Stephen A. Edwards
 * Columbia University
 */

module vga_framebuffer(input logic        clk,
	        input logic 	   reset,
		input logic [31:0] writedata, // 8 bits / pixel so we get 4 pixels at a time.
		input logic 	   write,
		input 		   chipselect,
		input logic [15:0]  address,  // 18000 chunks of 4 pixels at a time
		output logic [7:0] VGA_R, VGA_G, VGA_B,
		output logic 	   VGA_CLK, VGA_HS, VGA_VS,
		                   VGA_BLANK_n,
		output logic 	   VGA_SYNC_n);

   logic [10:0]	   hcount;
   logic [9:0]     vcount, pixel_col;

   logic [7:0] 	   background_r, background_g, background_b;
	
   vga_counters counters(.clk50(clk), .*);

   logic [1215:0] framebuffer [479:0]; // 480 rows, each with 150 pixels * 8 bits / pixel, rounded up to the nearest chunk of 64. So each row gets 38 chunks of 32 bits

   assign pixel_col = hcount[10:1] - 10'd245;

   always_ff @(posedge clk) begin
        if (reset) begin
         // Reset memory and other signals as needed
	 background_r <= 8'h0;
         background_g <= 8'h0;
         background_b <= 8'h80;
	 // Set default value in framebuffer
	 for (int row = 0; row < 480; row++) begin
	    for (int pixel = 0; pixel < 150; pixel++)
		framebuffer[row][pixel * 8 +: 8] = pixel % 3;
	    for (int buffer_pixel = 150; buffer_pixel < 152; buffer_pixel++)
		 // Give a default value to silence warnings
		framebuffer[row][buffer_pixel * 8 +: 8] = 8'd0;
	 end
        end else begin
            if (chipselect && write) begin
                if (address < 16'd38) begin
		   // 38 chunks per row
	           framebuffer[0][address * 32 +: 32] = writedata[31:0];
		end
            end
        end
    end

   always_comb begin
      {VGA_R, VGA_G, VGA_B} = {8'h0, 8'h0, 8'h0};
      if (VGA_BLANK_n) begin
	if (hcount[10:1] >= 10'd245 && hcount[10:1] < 10'd395 && vcount[9:0] < 10'd480) begin
	   // We are inside the 150 x 480 region of interest. Map the 8-bit value to a color
	    case (framebuffer[vcount[9:0]][pixel_col * 8 +: 8])
               8'd00: {VGA_R, VGA_G, VGA_B} = 24'hff0000; // Option 1
               8'd01: {VGA_R, VGA_G, VGA_B} = 24'h00ff00; // Option 2
	       8'd02: {VGA_R, VGA_G, VGA_B} = 24'h0000ff; // Option 3
               default: {VGA_R, VGA_G, VGA_B} = 24'hffffff; // Default to white
            endcase
	end else begin 
	   {VGA_R, VGA_G, VGA_B} = {background_r, background_g, background_b};
        end	
      end
   end
	       
endmodule

module vga_counters(
 input logic 	     clk50, reset,
 output logic [10:0] hcount,  // hcount[10:1] is pixel column
 output logic [9:0]  vcount,  // vcount[9:0] is pixel row
 output logic 	     VGA_CLK, VGA_HS, VGA_VS, VGA_BLANK_n, VGA_SYNC_n);

/*
 * 640 X 480 VGA timing for a 50 MHz clock: one pixel every other cycle
 * 
 * HCOUNT 1599 0             1279       1599 0
 *             _______________              ________
 * ___________|    Video      |____________|  Video
 * 
 * 
 * |SYNC| BP |<-- HACTIVE -->|FP|SYNC| BP |<-- HACTIVE
 *       _______________________      _____________
 * |____|       VGA_HS          |____|
 */
   // Parameters for hcount
   parameter HACTIVE      = 11'd 1280,
             HFRONT_PORCH = 11'd 32,
             HSYNC        = 11'd 192,
             HBACK_PORCH  = 11'd 96,   
             HTOTAL       = HACTIVE + HFRONT_PORCH + HSYNC +
                            HBACK_PORCH; // 1600
   
   // Parameters for vcount
   parameter VACTIVE      = 10'd 480,
             VFRONT_PORCH = 10'd 10,
             VSYNC        = 10'd 2,
             VBACK_PORCH  = 10'd 33,
             VTOTAL       = VACTIVE + VFRONT_PORCH + VSYNC +
                            VBACK_PORCH; // 525

   logic endOfLine;
   
   always_ff @(posedge clk50 or posedge reset)
     if (reset)          hcount <= 0;
     else if (endOfLine) hcount <= 0;
     else  	         hcount <= hcount + 11'd 1;

   assign endOfLine = hcount == HTOTAL - 1;
       
   logic endOfField;
   
   always_ff @(posedge clk50 or posedge reset)
     if (reset)          vcount <= 0;
     else if (endOfLine)
       if (endOfField)   vcount <= 0;
       else              vcount <= vcount + 10'd 1;

   assign endOfField = vcount == VTOTAL - 1;

   // Horizontal sync: from 0x520 to 0x5DF (0x57F)
   // 101 0010 0000 to 101 1101 1111
   assign VGA_HS = !( (hcount[10:8] == 3'b101) &
		      !(hcount[7:5] == 3'b111));
   assign VGA_VS = !( vcount[9:1] == (VACTIVE + VFRONT_PORCH) / 2);

   assign VGA_SYNC_n = 1'b0; // For putting sync on the green signal; unused
   
   // Horizontal active: 0 to 1279     Vertical active: 0 to 479
   // 101 0000 0000  1280	       01 1110 0000  480
   // 110 0011 1111  1599	       10 0000 1100  524
   assign VGA_BLANK_n = !( hcount[10] & (hcount[9] | hcount[8]) ) &
			!( vcount[9] | (vcount[8:5] == 4'b1111) );

   /* VGA_CLK is 25 MHz
    *             __    __    __
    * clk50    __|  |__|  |__|
    *        
    *             _____       __
    * hcount[0]__|     |_____|
    */
   assign VGA_CLK = hcount[0]; // 25 MHz clock: rising edge sensitive
   
endmodule
